module ConditionCheck(
  input[3:0] cond, statusReg,
  output hasCondition
);

  assign hasCondition = 1'b1;

endmodule
