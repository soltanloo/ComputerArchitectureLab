module ControlUnit(
  input s,
  input[1:0] mode,
  input[3:0] opCode,
  output WB_EN, MEM_R_EN, MEM_W_EN, EXE_CMD, B, S, Imm
);

  always @(*) begin
    
  end

endmodule