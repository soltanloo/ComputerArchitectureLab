module Val2Generate(
    input memrw,
    input[31:0] Val_Rm,
    input[23:0] Imm,
    input[11:0] Shift_operand,
    output[31:0] out
);


endmodule