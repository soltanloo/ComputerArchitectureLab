module ConditionCheck(
  input[3:0] cond, statusReg,
  output
);

